VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO CF_SRAM_4096x32
  CLASS BLOCK ;
  FOREIGN CF_SRAM_4096x32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 725.000 BY 925.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 21.400 10.640 23.160 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 21.400 438.010 23.160 479.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 21.400 888.010 23.160 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 71.400 10.640 73.160 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 71.400 438.010 73.160 479.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 71.400 888.010 73.160 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 121.400 10.640 123.160 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 121.400 438.010 123.160 479.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 121.400 888.010 123.160 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 171.400 10.640 173.160 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 171.400 438.010 173.160 479.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 171.400 888.010 173.160 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 221.400 10.640 223.160 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 221.400 438.010 223.160 479.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 221.400 888.010 223.160 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 271.400 10.640 273.160 29.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 271.400 438.150 273.160 479.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 271.400 888.150 273.160 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 321.400 10.640 323.160 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 321.400 438.010 323.160 479.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 321.400 888.010 323.160 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 371.400 10.640 373.160 29.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 371.400 438.150 373.160 479.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 371.400 888.150 373.160 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 421.400 10.640 423.160 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 421.400 438.010 423.160 479.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 421.400 888.010 423.160 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 471.400 10.640 473.160 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 471.400 438.010 473.160 479.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 471.400 888.010 473.160 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 521.400 10.640 523.160 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 521.400 438.010 523.160 479.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 521.400 888.010 523.160 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 571.400 10.640 573.160 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 571.400 438.010 573.160 479.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 571.400 888.010 573.160 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 621.400 10.640 623.160 29.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 621.400 438.150 623.160 479.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 621.400 888.150 623.160 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 671.400 10.640 673.160 29.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 671.400 438.150 673.160 479.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 671.400 888.150 673.160 914.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 26.760 719.680 28.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 76.760 719.680 78.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 126.760 719.680 128.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 176.760 719.680 178.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 276.760 719.680 278.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 326.760 719.680 328.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 376.760 719.680 378.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 426.760 719.680 428.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 476.760 719.680 478.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 526.760 719.680 528.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 576.760 719.680 578.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 626.760 719.680 628.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 726.760 719.680 728.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 776.760 719.680 778.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 826.760 719.680 828.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 876.760 719.680 878.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.990 226.760 359.800 228.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.990 676.760 359.800 678.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 684.990 226.760 719.680 228.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 684.990 676.760 719.680 678.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 23.970 0.000 27.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.970 0.000 57.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 83.970 0.000 87.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 113.970 0.000 117.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 143.970 0.000 147.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 173.970 0.000 177.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 203.970 0.000 207.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.970 0.000 237.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 263.970 0.000 267.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 293.970 0.000 297.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 323.970 0.000 327.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 353.970 0.000 357.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 383.970 0.000 387.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 413.970 0.000 417.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 443.970 0.000 447.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 473.970 0.000 477.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 503.970 0.000 507.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 533.970 0.000 537.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.970 0.000 567.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 593.970 0.000 597.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 623.970 0.000 627.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 653.970 0.000 657.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 683.970 0.000 687.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 713.970 0.000 717.070 925.000 ;
    END
    PORT
      LAYER met2 ;
        RECT 348.490 26.960 350.250 440.880 ;
    END
    PORT
      LAYER met2 ;
        RECT 702.230 478.480 703.990 892.400 ;
    END
    PORT
      LAYER met2 ;
        RECT 348.490 475.760 350.250 892.400 ;
    END
    PORT
      LAYER met2 ;
        RECT 702.230 26.960 703.990 440.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 906.580 711.400 908.340 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 9.640 10.640 11.400 29.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.640 438.150 11.400 479.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.640 888.150 11.400 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 59.640 10.640 61.400 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 59.640 438.010 61.400 479.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 59.640 888.010 61.400 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 109.640 10.640 111.400 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 109.640 438.010 111.400 479.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 109.640 888.010 111.400 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 159.640 10.640 161.400 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 159.640 438.010 161.400 479.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 159.640 888.010 161.400 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 209.640 10.640 211.400 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 209.640 438.010 211.400 479.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 209.640 888.010 211.400 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 259.640 10.640 261.400 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 259.640 438.010 261.400 479.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 259.640 888.010 261.400 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 309.640 10.640 311.400 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 309.640 438.010 311.400 479.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 309.640 888.010 311.400 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 359.640 10.640 361.400 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 359.640 438.010 361.400 479.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 359.640 888.010 361.400 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 409.640 10.640 411.400 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 409.640 438.010 411.400 479.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 409.640 888.010 411.400 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 459.640 10.640 461.400 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 459.640 438.010 461.400 479.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 459.640 888.010 461.400 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 509.640 10.640 511.400 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 509.640 438.010 511.400 479.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 509.640 888.010 511.400 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 559.640 10.640 561.400 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 559.640 438.010 561.400 479.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 559.640 888.010 561.400 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 609.640 10.640 611.400 29.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 609.640 438.150 611.400 479.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 609.640 888.150 611.400 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 659.640 10.640 661.400 29.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 659.640 438.010 661.400 479.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 659.640 888.010 661.400 914.160 ;
    END
    PORT
      LAYER met2 ;
        RECT 709.640 10.640 711.400 914.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 15.000 719.680 16.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 65.000 719.680 66.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 115.000 719.680 116.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 165.000 719.680 166.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 215.000 719.680 216.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 265.000 719.680 266.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 315.000 719.680 316.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 365.000 719.680 366.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 415.000 719.680 416.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 465.000 719.680 466.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 515.000 719.680 516.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 565.000 719.680 566.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 615.000 719.680 616.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 665.000 719.680 666.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 715.000 719.680 716.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 765.000 719.680 766.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 815.000 719.680 816.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 865.000 719.680 866.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.970 0.000 12.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.970 0.000 42.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 68.970 0.000 72.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.970 0.000 102.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 128.970 0.000 132.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 158.970 0.000 162.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 0.000 192.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 218.970 0.000 222.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.970 0.000 252.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 0.000 282.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 308.970 0.000 312.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 338.970 0.000 342.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 0.000 372.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 398.970 0.000 402.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 428.970 0.000 432.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 0.000 462.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 488.970 0.000 492.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 518.970 0.000 522.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 0.000 552.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 578.970 0.000 582.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 608.970 0.000 612.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 0.000 642.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 668.970 0.000 672.070 925.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 698.970 0.000 702.070 925.000 ;
    END
    PORT
      LAYER met2 ;
        RECT 336.530 26.960 338.290 440.880 ;
    END
    PORT
      LAYER met2 ;
        RECT 336.530 475.760 338.290 892.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 894.340 711.400 896.100 ;
    END
  END VPWR
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 396.610 0.000 396.890 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 410.410 0.000 410.690 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 424.210 0.000 424.490 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.810 0.000 452.090 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 0.000 465.890 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.410 0.000 479.690 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.210 0.000 493.490 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.010 0.000 507.290 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.810 0.000 521.090 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.410 0.000 548.690 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.210 0.000 562.490 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 0.000 576.290 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.810 0.000 590.090 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.610 0.000 603.890 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 0.000 617.690 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 0.000 631.490 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.010 0.000 645.290 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.810 0.000 659.090 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.610 0.000 672.890 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.410 0.000 686.690 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 327.610 0.000 327.890 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 355.210 0.000 355.490 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 369.010 0.000 369.290 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 401.210 0.000 401.490 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 415.010 0.000 415.290 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 428.810 0.000 429.090 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 442.610 0.000 442.890 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 456.410 0.000 456.690 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 484.010 0.000 484.290 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 497.810 0.000 498.090 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 511.610 0.000 511.890 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 525.410 0.000 525.690 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 263.210 0.000 263.490 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 539.210 0.000 539.490 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 553.010 0.000 553.290 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 580.610 0.000 580.890 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 594.410 0.000 594.690 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 608.210 0.000 608.490 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 622.010 0.000 622.290 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 635.810 0.000 636.090 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 649.610 0.000 649.890 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 663.410 0.000 663.690 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 281.610 0.000 281.890 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 677.210 0.000 677.490 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 691.010 0.000 691.290 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 300.010 0.000 300.290 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 346.010 0.000 346.290 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 359.810 0.000 360.090 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 387.410 0.000 387.690 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 419.610 0.000 419.890 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 433.410 0.000 433.690 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 447.210 0.000 447.490 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 461.010 0.000 461.290 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 474.810 0.000 475.090 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 488.610 0.000 488.890 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 516.210 0.000 516.490 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 530.010 0.000 530.290 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 543.810 0.000 544.090 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 557.610 0.000 557.890 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 571.410 0.000 571.690 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 585.210 0.000 585.490 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 612.810 0.000 613.090 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 626.610 0.000 626.890 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 640.410 0.000 640.690 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 654.210 0.000 654.490 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 668.010 0.000 668.290 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 286.210 0.000 286.490 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 681.810 0.000 682.090 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 304.610 0.000 304.890 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 336.810 0.000 337.090 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 350.610 0.000 350.890 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 290.810 0.000 291.090 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 719.440 914.005 ;
      LAYER met1 ;
        RECT 5.520 4.800 719.440 914.160 ;
      LAYER met2 ;
        RECT 11.680 887.870 21.120 891.470 ;
        RECT 10.100 887.730 21.120 887.870 ;
        RECT 23.440 887.730 59.360 891.470 ;
        RECT 61.680 887.730 71.120 891.470 ;
        RECT 73.440 887.730 109.360 891.470 ;
        RECT 111.680 887.730 121.120 891.470 ;
        RECT 123.440 887.730 159.360 891.470 ;
        RECT 161.680 887.730 171.120 891.470 ;
        RECT 173.440 887.730 209.360 891.470 ;
        RECT 211.680 887.730 221.120 891.470 ;
        RECT 223.440 887.730 259.360 891.470 ;
        RECT 261.680 887.870 271.120 891.470 ;
        RECT 273.440 887.870 309.360 891.470 ;
        RECT 261.680 887.730 309.360 887.870 ;
        RECT 311.680 887.730 321.120 891.470 ;
        RECT 323.440 887.730 336.250 891.470 ;
        RECT 10.100 480.140 336.250 887.730 ;
        RECT 10.100 480.000 21.120 480.140 ;
        RECT 11.680 437.870 21.120 480.000 ;
        RECT 10.100 437.730 21.120 437.870 ;
        RECT 23.440 437.730 59.360 480.140 ;
        RECT 61.680 437.730 71.120 480.140 ;
        RECT 73.440 437.730 109.360 480.140 ;
        RECT 111.680 437.730 121.120 480.140 ;
        RECT 123.440 437.730 159.360 480.140 ;
        RECT 161.680 437.730 171.120 480.140 ;
        RECT 173.440 437.730 209.360 480.140 ;
        RECT 211.680 437.730 221.120 480.140 ;
        RECT 223.440 437.730 259.360 480.140 ;
        RECT 261.680 480.000 309.360 480.140 ;
        RECT 261.680 437.870 271.120 480.000 ;
        RECT 273.440 437.870 309.360 480.000 ;
        RECT 261.680 437.730 309.360 437.870 ;
        RECT 311.680 437.730 321.120 480.140 ;
        RECT 323.440 475.480 336.250 480.140 ;
        RECT 338.570 475.480 348.210 891.470 ;
        RECT 350.530 887.730 359.360 891.470 ;
        RECT 361.680 887.870 371.120 891.470 ;
        RECT 373.440 887.870 409.360 891.470 ;
        RECT 361.680 887.730 409.360 887.870 ;
        RECT 411.680 887.730 421.120 891.470 ;
        RECT 423.440 887.730 459.360 891.470 ;
        RECT 461.680 887.730 471.120 891.470 ;
        RECT 473.440 887.730 509.360 891.470 ;
        RECT 511.680 887.730 521.120 891.470 ;
        RECT 523.440 887.730 559.360 891.470 ;
        RECT 561.680 887.730 571.120 891.470 ;
        RECT 573.440 887.870 609.360 891.470 ;
        RECT 611.680 887.870 621.120 891.470 ;
        RECT 623.440 887.870 659.360 891.470 ;
        RECT 573.440 887.730 659.360 887.870 ;
        RECT 661.680 887.870 671.120 891.470 ;
        RECT 673.440 887.870 701.950 891.470 ;
        RECT 661.680 887.730 701.950 887.870 ;
        RECT 350.530 480.140 701.950 887.730 ;
        RECT 350.530 475.480 359.360 480.140 ;
        RECT 323.440 441.160 359.360 475.480 ;
        RECT 323.440 437.730 336.250 441.160 ;
        RECT 10.100 30.140 336.250 437.730 ;
        RECT 10.100 30.000 21.120 30.140 ;
        RECT 11.680 10.360 21.120 30.000 ;
        RECT 23.440 10.360 59.360 30.140 ;
        RECT 61.680 10.360 71.120 30.140 ;
        RECT 73.440 10.360 109.360 30.140 ;
        RECT 111.680 10.360 121.120 30.140 ;
        RECT 123.440 10.360 159.360 30.140 ;
        RECT 161.680 10.360 171.120 30.140 ;
        RECT 173.440 10.360 209.360 30.140 ;
        RECT 211.680 10.360 221.120 30.140 ;
        RECT 223.440 10.360 259.360 30.140 ;
        RECT 261.680 30.000 309.360 30.140 ;
        RECT 261.680 10.360 271.120 30.000 ;
        RECT 273.440 10.360 309.360 30.000 ;
        RECT 311.680 10.360 321.120 30.140 ;
        RECT 323.440 26.680 336.250 30.140 ;
        RECT 338.570 26.680 348.210 441.160 ;
        RECT 350.530 437.730 359.360 441.160 ;
        RECT 361.680 480.000 409.360 480.140 ;
        RECT 361.680 437.870 371.120 480.000 ;
        RECT 373.440 437.870 409.360 480.000 ;
        RECT 361.680 437.730 409.360 437.870 ;
        RECT 411.680 437.730 421.120 480.140 ;
        RECT 423.440 437.730 459.360 480.140 ;
        RECT 461.680 437.730 471.120 480.140 ;
        RECT 473.440 437.730 509.360 480.140 ;
        RECT 511.680 437.730 521.120 480.140 ;
        RECT 523.440 437.730 559.360 480.140 ;
        RECT 561.680 437.730 571.120 480.140 ;
        RECT 573.440 480.000 659.360 480.140 ;
        RECT 573.440 437.870 609.360 480.000 ;
        RECT 611.680 437.870 621.120 480.000 ;
        RECT 623.440 437.870 659.360 480.000 ;
        RECT 573.440 437.730 659.360 437.870 ;
        RECT 661.680 480.000 701.950 480.140 ;
        RECT 661.680 437.870 671.120 480.000 ;
        RECT 673.440 478.200 701.950 480.000 ;
        RECT 704.270 478.200 709.360 891.470 ;
        RECT 673.440 441.160 709.360 478.200 ;
        RECT 673.440 437.870 701.950 441.160 ;
        RECT 661.680 437.730 701.950 437.870 ;
        RECT 350.530 30.140 701.950 437.730 ;
        RECT 350.530 26.680 359.360 30.140 ;
        RECT 323.440 10.360 359.360 26.680 ;
        RECT 361.680 30.000 409.360 30.140 ;
        RECT 361.680 10.360 371.120 30.000 ;
        RECT 373.440 10.360 409.360 30.000 ;
        RECT 411.680 10.360 421.120 30.140 ;
        RECT 423.440 10.360 459.360 30.140 ;
        RECT 461.680 10.360 471.120 30.140 ;
        RECT 473.440 10.360 509.360 30.140 ;
        RECT 511.680 10.360 521.120 30.140 ;
        RECT 523.440 10.360 559.360 30.140 ;
        RECT 561.680 10.360 571.120 30.140 ;
        RECT 573.440 30.000 659.360 30.140 ;
        RECT 573.440 10.360 609.360 30.000 ;
        RECT 611.680 10.360 621.120 30.000 ;
        RECT 623.440 10.360 659.360 30.000 ;
        RECT 661.680 30.000 701.950 30.140 ;
        RECT 661.680 10.360 671.120 30.000 ;
        RECT 673.440 26.680 701.950 30.000 ;
        RECT 704.270 26.680 709.360 441.160 ;
        RECT 673.440 10.360 709.360 26.680 ;
        RECT 711.680 10.360 717.500 891.470 ;
        RECT 10.100 4.280 717.500 10.360 ;
        RECT 10.100 3.670 212.330 4.280 ;
        RECT 213.170 3.670 216.930 4.280 ;
        RECT 217.770 3.670 221.530 4.280 ;
        RECT 222.370 3.670 226.130 4.280 ;
        RECT 226.970 3.670 230.730 4.280 ;
        RECT 231.570 3.670 235.330 4.280 ;
        RECT 236.170 3.670 239.930 4.280 ;
        RECT 240.770 3.670 244.530 4.280 ;
        RECT 245.370 3.670 249.130 4.280 ;
        RECT 249.970 3.670 253.730 4.280 ;
        RECT 254.570 3.670 258.330 4.280 ;
        RECT 259.170 3.670 262.930 4.280 ;
        RECT 263.770 3.670 267.530 4.280 ;
        RECT 268.370 3.670 272.130 4.280 ;
        RECT 272.970 3.670 276.730 4.280 ;
        RECT 277.570 3.670 281.330 4.280 ;
        RECT 282.170 3.670 285.930 4.280 ;
        RECT 286.770 3.670 290.530 4.280 ;
        RECT 291.370 3.670 295.130 4.280 ;
        RECT 295.970 3.670 299.730 4.280 ;
        RECT 300.570 3.670 304.330 4.280 ;
        RECT 305.170 3.670 308.930 4.280 ;
        RECT 309.770 3.670 313.530 4.280 ;
        RECT 314.370 3.670 318.130 4.280 ;
        RECT 318.970 3.670 322.730 4.280 ;
        RECT 323.570 3.670 327.330 4.280 ;
        RECT 328.170 3.670 331.930 4.280 ;
        RECT 332.770 3.670 336.530 4.280 ;
        RECT 337.370 3.670 341.130 4.280 ;
        RECT 341.970 3.670 345.730 4.280 ;
        RECT 346.570 3.670 350.330 4.280 ;
        RECT 351.170 3.670 354.930 4.280 ;
        RECT 355.770 3.670 359.530 4.280 ;
        RECT 360.370 3.670 364.130 4.280 ;
        RECT 364.970 3.670 368.730 4.280 ;
        RECT 369.570 3.670 373.330 4.280 ;
        RECT 374.170 3.670 377.930 4.280 ;
        RECT 378.770 3.670 382.530 4.280 ;
        RECT 383.370 3.670 387.130 4.280 ;
        RECT 387.970 3.670 391.730 4.280 ;
        RECT 392.570 3.670 396.330 4.280 ;
        RECT 397.170 3.670 400.930 4.280 ;
        RECT 401.770 3.670 405.530 4.280 ;
        RECT 406.370 3.670 410.130 4.280 ;
        RECT 410.970 3.670 414.730 4.280 ;
        RECT 415.570 3.670 419.330 4.280 ;
        RECT 420.170 3.670 423.930 4.280 ;
        RECT 424.770 3.670 428.530 4.280 ;
        RECT 429.370 3.670 433.130 4.280 ;
        RECT 433.970 3.670 437.730 4.280 ;
        RECT 438.570 3.670 442.330 4.280 ;
        RECT 443.170 3.670 446.930 4.280 ;
        RECT 447.770 3.670 451.530 4.280 ;
        RECT 452.370 3.670 456.130 4.280 ;
        RECT 456.970 3.670 460.730 4.280 ;
        RECT 461.570 3.670 465.330 4.280 ;
        RECT 466.170 3.670 469.930 4.280 ;
        RECT 470.770 3.670 474.530 4.280 ;
        RECT 475.370 3.670 479.130 4.280 ;
        RECT 479.970 3.670 483.730 4.280 ;
        RECT 484.570 3.670 488.330 4.280 ;
        RECT 489.170 3.670 492.930 4.280 ;
        RECT 493.770 3.670 497.530 4.280 ;
        RECT 498.370 3.670 502.130 4.280 ;
        RECT 502.970 3.670 506.730 4.280 ;
        RECT 507.570 3.670 511.330 4.280 ;
        RECT 512.170 3.670 515.930 4.280 ;
        RECT 516.770 3.670 520.530 4.280 ;
        RECT 521.370 3.670 525.130 4.280 ;
        RECT 525.970 3.670 529.730 4.280 ;
        RECT 530.570 3.670 534.330 4.280 ;
        RECT 535.170 3.670 538.930 4.280 ;
        RECT 539.770 3.670 543.530 4.280 ;
        RECT 544.370 3.670 548.130 4.280 ;
        RECT 548.970 3.670 552.730 4.280 ;
        RECT 553.570 3.670 557.330 4.280 ;
        RECT 558.170 3.670 561.930 4.280 ;
        RECT 562.770 3.670 566.530 4.280 ;
        RECT 567.370 3.670 571.130 4.280 ;
        RECT 571.970 3.670 575.730 4.280 ;
        RECT 576.570 3.670 580.330 4.280 ;
        RECT 581.170 3.670 584.930 4.280 ;
        RECT 585.770 3.670 589.530 4.280 ;
        RECT 590.370 3.670 594.130 4.280 ;
        RECT 594.970 3.670 598.730 4.280 ;
        RECT 599.570 3.670 603.330 4.280 ;
        RECT 604.170 3.670 607.930 4.280 ;
        RECT 608.770 3.670 612.530 4.280 ;
        RECT 613.370 3.670 617.130 4.280 ;
        RECT 617.970 3.670 621.730 4.280 ;
        RECT 622.570 3.670 626.330 4.280 ;
        RECT 627.170 3.670 630.930 4.280 ;
        RECT 631.770 3.670 635.530 4.280 ;
        RECT 636.370 3.670 640.130 4.280 ;
        RECT 640.970 3.670 644.730 4.280 ;
        RECT 645.570 3.670 649.330 4.280 ;
        RECT 650.170 3.670 653.930 4.280 ;
        RECT 654.770 3.670 658.530 4.280 ;
        RECT 659.370 3.670 663.130 4.280 ;
        RECT 663.970 3.670 667.730 4.280 ;
        RECT 668.570 3.670 672.330 4.280 ;
        RECT 673.170 3.670 676.930 4.280 ;
        RECT 677.770 3.670 681.530 4.280 ;
        RECT 682.370 3.670 686.130 4.280 ;
        RECT 686.970 3.670 690.730 4.280 ;
        RECT 691.570 3.670 695.330 4.280 ;
        RECT 696.170 3.670 717.500 4.280 ;
      LAYER met3 ;
        RECT 10.100 878.920 714.775 887.225 ;
        RECT 10.100 867.160 714.775 876.360 ;
        RECT 10.100 828.920 714.775 864.600 ;
        RECT 10.100 817.160 714.775 826.360 ;
        RECT 10.100 778.920 714.775 814.600 ;
        RECT 10.100 767.160 714.775 776.360 ;
        RECT 10.100 728.920 714.775 764.600 ;
        RECT 10.100 717.160 714.775 726.360 ;
        RECT 10.100 678.920 714.775 714.600 ;
        RECT 10.100 676.360 324.590 678.920 ;
        RECT 360.200 676.360 684.590 678.920 ;
        RECT 10.100 667.160 714.775 676.360 ;
        RECT 10.100 628.920 714.775 664.600 ;
        RECT 10.100 617.160 714.775 626.360 ;
        RECT 10.100 578.920 714.775 614.600 ;
        RECT 10.100 567.160 714.775 576.360 ;
        RECT 10.100 528.920 714.775 564.600 ;
        RECT 10.100 517.160 714.775 526.360 ;
        RECT 10.100 478.920 714.775 514.600 ;
        RECT 10.100 467.160 714.775 476.360 ;
        RECT 10.100 428.920 714.775 464.600 ;
        RECT 10.100 417.160 714.775 426.360 ;
        RECT 10.100 378.920 714.775 414.600 ;
        RECT 10.100 367.160 714.775 376.360 ;
        RECT 10.100 328.920 714.775 364.600 ;
        RECT 10.100 317.160 714.775 326.360 ;
        RECT 10.100 278.920 714.775 314.600 ;
        RECT 10.100 267.160 714.775 276.360 ;
        RECT 10.100 228.920 714.775 264.600 ;
        RECT 10.100 226.360 324.590 228.920 ;
        RECT 360.200 226.360 684.590 228.920 ;
        RECT 10.100 217.160 714.775 226.360 ;
        RECT 10.100 178.920 714.775 214.600 ;
        RECT 10.100 167.160 714.775 176.360 ;
        RECT 10.100 128.920 714.775 164.600 ;
        RECT 10.100 117.160 714.775 126.360 ;
        RECT 10.100 78.920 714.775 114.600 ;
        RECT 10.100 67.160 714.775 76.360 ;
        RECT 10.100 28.920 714.775 64.600 ;
        RECT 10.100 17.160 714.775 26.360 ;
        RECT 10.100 11.055 714.775 14.600 ;
      LAYER met4 ;
        RECT 314.935 11.735 323.570 798.145 ;
        RECT 327.470 11.735 338.570 798.145 ;
        RECT 342.470 11.735 353.570 798.145 ;
        RECT 357.470 11.735 368.570 798.145 ;
        RECT 372.470 11.735 383.570 798.145 ;
        RECT 387.470 11.735 398.570 798.145 ;
        RECT 402.470 11.735 413.570 798.145 ;
        RECT 417.470 11.735 428.570 798.145 ;
        RECT 432.470 11.735 443.570 798.145 ;
        RECT 447.470 11.735 458.570 798.145 ;
        RECT 462.470 11.735 473.570 798.145 ;
        RECT 477.470 11.735 488.570 798.145 ;
        RECT 492.470 11.735 503.570 798.145 ;
        RECT 507.470 11.735 518.570 798.145 ;
        RECT 522.470 11.735 533.570 798.145 ;
        RECT 537.470 11.735 548.570 798.145 ;
        RECT 552.470 11.735 563.570 798.145 ;
        RECT 567.470 11.735 578.570 798.145 ;
        RECT 582.470 11.735 593.570 798.145 ;
        RECT 597.470 11.735 608.570 798.145 ;
        RECT 612.470 11.735 623.570 798.145 ;
        RECT 627.470 11.735 638.570 798.145 ;
        RECT 642.470 11.735 653.570 798.145 ;
        RECT 657.470 11.735 668.570 798.145 ;
        RECT 672.470 11.735 683.570 798.145 ;
        RECT 687.470 11.735 698.570 798.145 ;
        RECT 702.470 11.735 706.265 798.145 ;
      LAYER met5 ;
        RECT 318.900 24.700 697.700 441.100 ;
  END
END CF_SRAM_4096x32
END LIBRARY

